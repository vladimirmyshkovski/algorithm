module main

fn test_new_user() {}
