module main

fn test_new_product() {
	first_product := Product{
		product_hashes: []
		work: Work{
			signature: 'fake_signature'
			hours: 10
		}
		purpose: ProductPurpose.consume
		class: ProductClass.b
	}
}
